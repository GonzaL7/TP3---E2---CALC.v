module memory (



)

endmodule;