module testbenchALL;

endmodule